//-----------------------------------------------------
// File Name   : alucodes.sv
// Function    : pMIPS ALU funcRon code definiRons 
// Version: 1,  only 2 funcs
// Author:  ks6n19
// Last rev.  11/05/20
//-----------------------------------------------------


`define RADD  1'b0
`define RMUL 1'b1
